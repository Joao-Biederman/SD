entity nome is
	port(
		c0 : in bit;
		z : out bit
	);
end entity;

architecture nomeComportamento of nome is
begin

end architecture;